PK   Z�S$��`�=  �u    cirkitFile.json��r$���_EF��U��9���ս3���L��\��hq�hSMֲX����@�2�L���)32"��?�-�uQF�デ�� <�rq��i���o�ƫ?�w�oo.�"���������O����7W��W�k?��⫿�����0��nl���\�)h������(?Dݦ�L1tW�J_|���}�K�W$f�J�W�%<��p���Nݵ���_}�}��]��7�x!�wǊU*�����A*A_���������f���ғ�����r�Z�6nR����䧩�J��=8�.QTz�A9�j;U����)�|�Fh^�� ~R	�*��4?ȗVp��v(�A��kQ*�ݴ|�؉�|7�<�ٛ����="�ah�a<�'�iی�Q��:K�jb��թ��h0y�v_:��^��'N�|��`
'4+-5+��I�ه�"�B>��E0E>O�	�H�I��">;�2$��IP,���bc0���S.�4u����q�s�XS�����gZ�I�&�R�|��`
�l#���D��Lҧ)�j�"�B>]�E�++O���<M�д�B,�)��^,�) �jV4mJS>+�*�"�B���"�B���"�B���"�B��"�B��"����l����]����]����]�� �А�N'��bL!��bL!��bL!��bL!��b���}�XS�}�XS�}�XS�}�XS�}�XS�}�XS�}�XS�}�XS�}�XS�}�X��
r�)�r�)�r߹&��=��R��@	��ު�WOB	�{�
�{�b�;���ȭbe6,d�J���|�uA
���\���i��R	��U�~��An�b�Ѭn�*�T�^�vU� ��߸%
M�V���� �I��"f[�>ür��|V\�}UJ!��ֶ;�Rȧ��S�[t���,�h(Ձ|J�x�q%g:��qVf����͊���٦���jRG�mP�`H�f�[r�ib:��'"�������tR�v��H�uRD�O��u��LOP:���N����A��g}��Ch�b��bu�#,'�X�9��t����;�����t�*`u������`]���~|Κ�LUоѼo2U%���j�t���WVwVwP:���バ�|�rCi(����$��-�	Յ΋f��l]�lt^N���Z"��'<���y�ne�yx�������|y��?p���#0_^����a��ߩ�Ģc��Y���	�m��ϻ�ٚF�@8�$hF`>��3�`��E,���y����"���|��.V�.b��w���?h�GҔ�=:�=���	��}a� V?�m8e3��̀S6,��rY���)���|��X���G`�\�?��5,��r!�������|��
X���G`�\ �?p���#0_.]��~�|�˕s��o���/������G`�\��?�>�>p�a����X>��*O`���,��r}*�������|��X���G`�\�?p���#0_�f�8����/�a��ρ�,��r9�������|��X���G`�\��?p���#0_�7��P�T8�p��Á�,��r�G�������|�:%X���G`�\W�?p���#0_�
�8����/�2��σ�,��rV�������|�~,X���G`�\��?p���#0_���8����/W�]� ]� �xp�������|��3X���G`�\��?p���#0_���8����	�gi�d��ϵı����G`�\�?p��#0_��~�'�[�H���x��ؤ&�=��D�m�S۱��>`-p��B���s�n�*�RP+�F����.<ϲO$6�[/}�3���؋:�$�>��̙͏��������͏��;�DW5Q4�e���{ѽ��ޢ�M'��l�YѽeŬ��i���W�?�Ѳ��u��l~\p��:ӲǠK���:�0�=,�E͗瀢�Io%��/d˂�4$�H��7$�m/���AQ��%\v륹���K�P٭�㍄�d#��#���K��bP6��>�+u�nO���R�_�y���:��ޕ�o�{��;�ݒ�)��%��{ˬ=��-�\M��[fj��֢f�!�])
�m#[,���m#Y���H����8G��.���8Gr�1���'��.�ʍS���t��1�����]IR��/�q���lCj�S.Y��NY���P�zcV�^�|��\��S����U;���[��?^�{Q�廇IS�"�h#7o������u!�8�i�k�E�W�E�'�n�XQ�j�fT���'c�[�{Q�S�4ʅ��k�j�1p_�4Nf����^�|����ɵ�o�1��&n�S��abC�~�[�����w}[?������;�-7�8$3��Kk�/j����Swf�����m;���]c�f�M��(U�|���}���V���-m�./�q���Z�r����wg�ZO[iJl6�s�h�ǆ&4�vkVW�|���`�4E��d9�-?8�@T�G�L;%=u+w/j�rw��qh&n޲��,��Dm?6��Zߋ�/�=��b0�r���2����ώ#Nkw/j�2�D4�:;����U"�f����ݽ�����1���^c����hy��iBkmy�4�=��݋�����5=畊��st��lZ�:���6d��fuE͗�>L��{���!�s��y�1c�M\g�C�*h�bu���8�Lm���Q��C�xz�4�0�Y]Is�ݗ�Ѣ��k~���uש�Xn�BT�p�֏��M�<��⺢�+�{I��5_8oh�V���S����7�	z�hy��5_�{Q��5_�{�΍���v���j=��}m�k;�|]I�O[�|��E͗���^��yV2�9��9$�	z�Ym�e�1�6�K������+㽤�r��ۮ���D�i����簐z�G��b7�����+�LI��5_�&�m��Dˡ'<E��5>m4�#����|u�o7������W��W���ۻ���"y�������z�u��ed����)H�n���Ͽ�^NdPD�#���V+H�n����hht2"�"
(��6{a�@�v���X�9�%Q��H�~��E>H�^̴��%��7�	������L K��S��m� 1�|7�}.i��	�	�u	&i�������wZ'鸃�p�^z�9��F4��̏�����}��p�3�����､��:|/�L���b�E���Q��n?�i')F�1̏�$���̏X(���v1!̏�$��F̏[X<����ѯ�	��Q�r�~n%��� �q�"d��q��\������Q�rYq,�0?����_Ø`~���8JR.�c��q��(I��0�	�&�[��q��(I��,�	��̏�$咧0&�w0?���Ks��P�r�K̏{�GI�eaL0?�a~%)��1�����q��\������Q�r96̏�GIʥ�`L0?`~�@R�����+�"A%��J�P�T�����l�|/$�=��)��$�a_�궂B"�����h{�,$	z�W$�#���}E�D A�`;P!H�þ���i�D��m���Z�I�O����M0�]����	�v�2�|�~7��ޔR&��S��	�Q���l|A����W�v��O�CXg� ��j\ �W�=eA"�O�r�`�*�KW�����Y�R�z=��	\*P�5X�
+�5U�z���j�RV�Ϊ���[(�`�*��cV���7R0��JUX9S����o�`��t�U��㯩���+Ua�W�_Y�K�+Ua�k/u�SY�\Uh�4- 窔t��d�^�
-��(�F2s(��i"��(�N�Eu��*�T�6�M��m��
-ա�_�A�NV�v�)!�\V'�S����i!��N.Fu�1���PZ�C����m���
-ա�g���NVV�����3�Utk��eUh�m>k^G�u�*�t���:y����U��Ӵ %���L���
-ա�5��N^V�����Zut['/�BKuhsM�:���
-ա͵1��N^V�����ut['/�BKuhs��:����U��:���J��Iu�*�T�6׎���:���R�\��n��T�BKuhs-�:���[��v�:y�����:yYZ�C�k+��m���
-ա�5���N^V�����ZWut['/�BKuhsͮ:����U��:���X���˪�R�\C��n]���
-ա͵���N^V�����vut['/�BKuhsm�:����U��:���`�V:IV�(Y������\���
-ա�5��N^V�����ڕut['/�BKuhs�:����U��:���h���˪�R�\��n}���
-ա͵]��N^V������ut['/�BKuhs��:����U��:��fp���˪�R�\���n+U��T�N^���e�N^V�����Z�ut['/�BKuhsM�:����U��:��6x���˪��iZ�y�P'/u�*�T�6�j���:yYZ�C�k��hC��eUh���������xse:m�14��&*giRMLQ�:����p�T
���R���L)�z�ߚ�m�@����fo���V e��$gJY�m~���z�gJY�!~������/�w1��k�_H���7$���D�×���J����o����Y���,FO�:�
.L�QkU۸I�&Nn���~�gJY��~����gJY�Z~���7��x�3��2ER6�L�������L);/3���V2^��.��?W�~��w����Y�7��6ȞƄ	cô3���������/d^O�]�������L�Ί�w���y���W�+�nMreb6��21~+ (�21q+8*��B�21�VT^6�b|��7��ئ���jRG�mP�`H�f�[r��P�Jo��ER�8s���i�H��r�ERܖ7wf�ƓWS�F��)r�t��1�����ݎ��l>�V��ن��'�\�Z%��읦�:���R$e�e�K�w��c���Jcg�5�E��?�f)���&M�����,�m���`ׅd⠧���ER�G#۾O^�N�.Ռͨ��O�O�W�R$e[/G=��r!u��[��v�A3��ll���H�dq^O��A��θib)��)&����1��qT"e�e�ml�D�z�[����ApqHfS�
�Q���Hz�������=�ж����1}3Ŧ-�IK�l�����k��Z�Rly��;�'�����,ER6Y���S�&�[q�?�AEvݡ	M�]��I�d�ۧ):�&�I����mT�G�L;%=u�,ER�Y�nơ�XJ��۳(�QT6��ؐKz)��ɒ�av10������eοg��")�scdj�ڵShy&��J���Z������")�,���Dl������hy��Y�X��e���R$e��ہC�)�d&��֨���=�n��M�a"?��+� y4��v�'��{��Y����l�.ux��a�M�kT;��h��y�:��["ò5I�\K	nԬ�NƲ����c�~to��Z�Iَ_J�l�Hʦ^�dx�[5R�R�T�ު�t&���9�Hʦ^��l�Hʦ^Z�tnd�����T�9���h{?X��X�wK�l�%R6�R$eS/i�5���T���@��	�<��5�[�;���3�l��)���Dʦ^�ۮ���ι<�qD6�5So��8���D���X"eS/ERJ��	c���rt�9��-���C�� �ȿlK)�/�R^��;1W��W����⫿<�}����7�����K�sJ�~� �$h�� B��� !	����X@�@���5 D A��"���>H�~O
�$�a�E�6�m��6�7J�޿`�0�|7��7J��>%�́�$���̇̉�$��v	̏�GI���&\���a~���8J���W�0�����q�$��I�a��q��(Iz�������Q��~�&��q��(I�:8�	���[J��q��(I��3�	��-̏�$��0&��0?�����`~���8JR��
c��q��(I�
'�	�&�[��q��(I�Z"�	��̏�$��|0&�w0?������^������q��\}�����Q�r�+��&��&̏{�GI�U�`L0?�a~%)W��1��x��q��\u�����$��K��h�;��j;U����)�E�����+*$�Vw!HPɾ�B"�S۞2�@�J����+*$	*�WTHT����$�d_Q!HPɾ�B"���}E�.�qn�v�2�<w�n�R&��.�T�����J�`��`7P)ӂ��+��*,�����RV���Ϻ�^g�!��JUX9����YaE�j�RV���uV����T���*z���h�+Ua�쬊^gE�!��JUX9Ǭ��Y�{�j�RVΔ��uV����T����*z���h�+Ua�W���h�@��`�*�y�NbP'�BKuh�R�Vʺ*�]u�.��xQ�̫
-ա�kzut['��BKuh��d������Rڼ�ZG�u��*�T�6���m�L�
-ա�gi��N6V�����3�ut['#�BKuh���:����U��:���v�u�*�T�6�5���:yYZ�C�����m�7b�^����L�����˪�R�\à�n��eUh�m��PG�u�*�T�6ה���:yYZ�C�kc��m���
-ա�5>��N^V�����Z%ut['/�BKuhs͕:���eUh�m�SG�u�*�T�6�����:yYZ�C�k���m�݊��+���l�����˪�R�\[��n��eUh�m�UG�u�*�T�6׺���:yYZ�C�kv��m���
-ա͵���N^V�����jUt���eUh�m�WG�u�*�T�6״���:yYZ�C�k���m���
-ա�5���I�JG���e�N^���eUh�m��XG�u�*�T�6׮���:yYZ�C�kp��m���
-ա͵D��N^V����暨Ut���eUh�m��ZG�u�*�T�6ר���:yYZ�C�k���m���
-ա�5���N^V�������ut[��G�2u�2_'/�u�*�T�6ע���:yYZ�C�kj��m���
-ա͵���N^V������Ut��eUh�m��^G�u�*�T�6ל���:yYZ*��o�p{3��_�N�f�꼉�Y�TST�N}?$G�Y,����Z�gJY�N|���z�gJY� |�����gJY��{�����gJY�G~�����Z�x1ֻT\�\1�[*}��M�ӓ�����r�Z�6nR����䧩��2ER6�S����T$e��I�|�ER6u�̓��2ER6�L��M/Sfu ��Xﶗ)���mgU&c� gE&�ƊƊ�c��`��`��`��`��`��`��`�x���ٴb�tԵ�SM�H�����}Kn2*mG5ER0,��H��x*��9������ԥQ�q��6��q��'��`��[$eS��n����ON�d�J>8e�vSC���f)���2����;��QΌ^���j����i�o�I�d	���ER�F��6Iuw��B2q�����")�#��m�'�n�X��j�fT���'c�+`)�������A��:~ҭVM;��6�C�^J�l�8�'�ڠ�qg�4����a��\�8*���2�6�~"E��ܭ��I�� �8$3��KϨH�v2N]�Y]���hێ�|ט��b��%R6Y|���5Zu��	)�<z������}��m�")�,�B�c�O���8��"��Є&ڮ�v��l�t����J����[~��6*�#u�����m�")�,V7��L,�e��Y�(*��~lȥ�I�dI�0�{~҆G���߳��SK���12�a��)�<��^%rlu-���O�PK��M�~Lf"6�����t�<�򬦵�<�N}��Hʶ�[ӷ�S�9�Llu�QV2z,��")�,�D~�W:z�=G����?�ޤ�u֗D�ER�m�:<���ͦ�5��G���<L��-��aٌ���lF�����۩�X�²T�p�ڏ��M�<R��")��K��M�I�~3�D�V��������7�	z�D�d(����_"e{��Dʦ^Z�tnd�����T�9���h{?X��X�wK�l�%R6�R$eS/i�5���T���@��	�<��5�[�;���3�l��)���Dʦ^�ۮ���ι<�qD6�5So��8���D���X"eS/ERJ��	c���rt�9��-���C�� �ȿlK)�/�R^�������!���ۻ���?/���.�|}7~����������n�.������E�z?���[{�¤���dƢ{�*���Z��,�7ɖ��fu�������֝_���w���o��oۛ���|���w?����wڼ���8���}�8I�*��������$��UyE��<�%�h�|O`|��Hh���FE,�"6�^�k$��^��VHX��R�b;�a�V��8�lY�0��'V��F��RrkIxF��a�V&�(���f�H 3͂1|�Ds��)ɶ{JgYQ����o/����Q��5�����84%��uÿ���R�$Z;;(+YÑ�\�h���l�};�$��D �1��π���_�H�$������6H�@�!����̟A v�e��U�� ����`�(#���h�pf�а�p1D&�ы�1��#N��^�}����1�#�E�'�^)�ڎ�մ���i
��͗��J#K�_]ሣ���>��u��iH��G�#5�B�����x����a(���"�B��
���RLRj�bN4�ዙ��ǭ�w㏷���f8������z��~�wH7+�	��g ��C;��ߨa�B)|��a�)�>�'ك��_ H���T��o}P
w�.��/rw�h�}sJ�^�%�����u�X�Oz4|I��X��Ή�8�co!�[���-�i�q��3�
Æ{z�-�B���y�З�� �O�� �qdl���J�s.��
|�2wIO� Ԃ>�@B��0���1^E��S�׷�ٹ!9�����r�w?i'?�cLpD�i�U;�"���ҳMr�'9���<3G'�?u�����۟k���<LN =$pb���BL!=7���|�cJCr��FH�?�X�m�=��ɳXx��S�bg�A1��X(�Bx:��f�h���V_;hz����ϟ��g�?}ZO��aB�m�P	�J�-H
 ����wr�8@�S�p��s�[>P ���ȫ�`68a��lA���F^��G��6���U���g�o�} @����$L�������?�d��3�?Y.���g��U߂C�z*ԩ�P��� �N^���v��_v��*�@��vd�u��@���x P�<*tq��K��5z�� ��ꩻ�T^���JFyឺg���i� �_\�'������۟_���]���t}s{��/�z���4�=����է��⫿H�S�|�,s�л��
)�"��������7r(+W�XD�Z�b9�= �29�$
��\5b���)�"r�~��l�A%9T#W�XĮ����� �!�?2�:!��gP�)�eb�Rp^�p�r�j�EvA{�R,�w%��ݲ���)��h`�^�K�ci/�hpI�<�o�e�2��;Nj2@�lNxj�K4 O-��{#� �f���ܽ�.p�r:�V�s \���f��s�5�e�\�P���D��\���|�\s ��\��g��v������2��|�2v{�� �k�W.c�GP���m�2v�{�~�P�ܫ\�n����^���e춲�9 ����\�nG���O���e�6��9 ����\�nO��C.�9 �T.C�
r�?� *�� *�� *�� *�� *�� *�� *������e0���e䚕 �5�[��F�[{H���"ַ�oО�fi��
�֦�B
����#Ո���)�K/n
�&�B(������~-����I�[]ߏR%�Ww�R�E�7��d
-{m�,��b�J �7����?l@�b��*dll1)� x�S[L�^�om/~�^J	p�r;N��%:FC'E�i�C��	&>��������8��P9tL����#0��fe��7n��C�9��Ƀ�ӂ�т���#0'/`�9���|���
�?����|�����������;Dq=z����X\��
����L`s���O_5`�5`�a�̧*�`��Y: �����b<��deV0*��G>R�IJx
��a��:A�T��0Ѽ��y*�|���y�0!�	��Z���LHhB}�y\��	�p�E����b���}�*��G�S���9�>�|�Ѣ�"¦�&$4a>[��!:�0E���		M�g��
Ĭ��"0�aIG��2 ��=B�	`���q��������t�c�)�q5Zy��)�0�F���		M�O��u�Ny���&̧��:D���0��G��ŀ		M���u��b���&�%�:Dg1`BB���m*�,LHh�\��C��30!�	s��������&�5B�:��9�o:C�)��Xt�&$4a.Ƃ�!:O�0�A����		M���u��S���&�|�:D�)`BB��Ch��0!�	s�$�:O�0}B����		M�V�u��S���&�Ŷ�:D�)`BB�Bah����Ƞ���S:O�0hC����		M��ˡu��S���&̅��:D�)`BB�~h��0!�	sAB�=:O�0SD����		M�A�u��S���&�E,�:D�)`BB��h��0!�	s�P��g����y�G�)���		M����u��S���&�g�:D�)`BB�b�h��0!� <:&,�~����U�i��Є�f1Z��LHh�\o�����E���G��u��L�����7�����m�ШΛ���I51E����Cr4�SE�O�)n^���<��N|J\"���H n^xS���g����U�?���n��g�l?+�{�)�0m+�w¶%#�ć����;a�A"on�$-'*�҂}��[�U��I9j�j7)���C���ϋٟ�~V�������g��U>�����Nx�$��}�گx����)�vN�_�e�'6^��΋j�+@j�'�-��2y'�Ղ�+�'5��G��p%�NX�G/�'>� �ɛϰ���;>.D e����ҌX&�|�.�wKF����KO������"�2y��1�ɛ�����l��z��ǌ�ئ���jRG�mP�`H�f�[r���DvG�z���saR-�2�?1̽H܉�ha4:3D�ɫ�K�r�9�m:E�]O����ŧE�W�}���lCj�S.Y��NY�SC��Y�Q���O~pi�N5zl�3�Wi쬚�frM#�x��E�W�&��.��6r��I�k�;]����&���_{<<�>y5p��jT36�'?�>����گ��⨧qP.���_�Uӎ��c�q2�������+�w^O��A�ct7Mܞ@E���8�j�%�W�?�6�~"E��܉��M�F\��ԥU��_��ǩ�;������۶����1}3Ŧ]�OKگ�߷��]�U�j�<b��۳cv���C�֯ݿ�����E��S���q�?�AE���	M�ݪ��_�7�>Mѩ4��ϯ��m�B?Rg�)�[�Q���[݌C3q����g!���l j��!�V�_�~���Q��c������\v��{�$qZ�Q���'2�a��)��m�9���G��hh��E�W�ߏ�LĦ{��NG���9����Xv�k�/j���������}��OkT�S����q���گ�����JG�����<��ޛ4�����O�~�����;x��lD]�ڑGr;���k�a\�������D�E�W�7�5+�S��ܞ����H�ݛ`yl��E������+�/j��3���V����Z����7�	z��f���_�Q����_��΍��؈���j=O�}m�k;W�_I�5�[�~��E�W���^��y�2�9��9~��{�Yw�e2'>6{f���_�~m���_�b۵�S�9���_���G�G�ݴ��Kگ�?%�W�_�~}��0��-�O�M���r8��8���6��v����~�����xnw=\��^���_�����W���K�y(/-�媼����@^��+*y�rW�� �{��{-�[��p�û������=����w+>�u����n�w���[ݽ��}�m����K��7.v/�w����K�PN�s����ܠd��Aɒ�A��5��%I��
��%i�A��<��AI�yР$S<hP��4(��$OJ��C�+HO���O� 8hP�v� ĝ�l���Ɇ%A�Ɇ%��Ɇ%��Ɇ%��R7'�Æy5cr�&z|7&�N�}�h�f�}H��g�5;-��C��35�?ݤf������'�O���f��S�վ�ѻ������$�Dގ�y1�Iz&z�Ԝ�1��t��Jhh᱗�ߛ�8���j8��E8����N�^ƺ8q�pC�h�����%	��`���H��A
�e�P��g�|���q���|���S
_b��P�i�\J�;p��9͒G)�o zr[���<J��
��Ap�Q������n(�
�훆�DF�����D$%���X�)�d�*��I��a�+�
fE�9A�D���M�(��5��~�H?�P��qnE&
�$
;�/n=8�.��y�A���ִ���i
}��􉧯�����fO;��$%ԋ��g��'�s����	��ũ��P8���o0�g�B@��1��ۜpq�-kB7��'�B>�#�J[��<WH����K�s�ř��Pj��:¹F4_�Չ��J����z��O1%)��1���lNȟ�1�JލԞ��|��f�����_�o��}~ɠ�~]|u����g��GW���/��Kf~�>\��K�ᒛ_����Rx���å8��.�����R3�D��4��Gz���#>��鑟���м���w��@�>��'j��<>R3����*=^��5�33יyԙ9��'�:��O3קyԙ9��ǾӉ�?����i�i����2�\�}생��>���uf��\g�Qgv�3��;׋}�3;�3��3;י}ԋ���>�Ş�����_�״��_�pT�7�������F��r�Sޯ��W�ؒ�n��n�Wy�����>�Wd���;Q� ���8�3T�G}�mL�l^��+Θ��G�e�6������+N(��<&�����aA?K}xʚ>���ϻL���ѯ�n?�w��cޓ���)���������F��&wi����1:���ؘl�c�R�,�Aչ4��e���v��o>޷7��M��w�w׌��.>}Ȇs}׿:�{�g�����mC�����ҾTG|�`���߭��/��%9�\�������^���ㅘ.ͩ��/<���xx�ǟzꎷ�m$����ח����=����^��ǟ7��3{9?�4������4\���x�q�d�ԗĞ�}\���&���<�Ϗ�w�7y���1�;_}w�������3C�>���5����?���W7߲܋��l�|��x�o�������������nd;��q�V�c{�ij��Ow��������n�t}s 9 ʸt��j���_c��;�>����N�l�S�����s�xp�U,ʄ<:��f��7GF�x����z�b���Ԇ��6ۄ�6v�
IsOW�Y����ĥ~��ݍT���m��a�WLGJ�h�[ja�X�W(,]�Km(-�9�0��x��Sz�2J�W�O����)=\�?���/|��;�֤�F;��Ar|�ͺ�}�0���h��7O��[䭦������`'�F�f��hko�h�d._x#���}0�x����R��fn��I������h���-���l�1�݅�x�if��]2�%τ|���M�������I��	�.��ݶw>�4<��&>vx��(�<��`�If��R}�����B��4�1���K�L�hcx����ȣ��Iǳ�}����}�9w` <���I�� @���Q��l!GAIx3����y��@�~�HZr!��r�,e!ƺC��B�N�X�1.ĸC�Io��B�f"����]%r��G9J(җ��+�wkָ��ԩ���Ѫ��Vu�N�O������MS�3Rr��d����`o�8{�|�����zO�����>��ы�����n�������{�x�揟Į������,�~�h9O5�E����W���}?��0�p��g������)��CV��ݡ�K��w~���_����������b�	˚�/?�؍w?����oڛ��*���}�t�����j�3�)q�L�gk�7]:j�55�|t� �7�ݼ�k[��#�������ا޷�T��ti��y8���S�}��f��@VL��d�6�&��FH�6%�cJ�F'5�3�%���i���8!��ov�dǜ�>ϩ���{cc5[sp!�&I͸�$~��%w���u���,3޽�wA[���w�s^¥�>J��`�v\T �$u�w|�\������8rw�*|�	9؝?N�	�7�mِԎ�ꖔر���;w|�߼�?�[���<�+(&�v�1+�p��	^H☢��N�2�>^�ڻ��e��J��͈_͈UN��.J�W�n7��o<��t�Sc���qI����y#��,ni>s���|�}��׳��nQk������
��DQ��"㥼u�y����6א��������&V ��<�ņ=�fN)9���6Rk-*uWb��5�p�}G�7"���9�ܔ_�7ο��$6ޢ��E���=�q���k�]�ތ�ՌיKm8m�	16��$l�PT�d�7>��p��6���.����n����r]���d��ə�Vj�E�h,7�|<��{�]�����w����_�V�g���o/^�̷����ۧcs ����\��33��y����ɏ,g�q���0��X=��ǩk�~���T.������OZ<_�OW��o����>���r�(*.]bi���}<�����Ne=_z�Wzs U�@����;�+0/Ŀ���̣�yXsM���J���^��{a/]Ǜ�h9�c�x�"�H��
P�A����3��ŅƼ�Im3�E_~(7�}����l�������YN�����^���a]����^��_tY�{��w�h�OYz{i^,Gl��cz;8�����2n0��O�0����`��%�A>p�.��7Atj�Z�Mt���;>���L�g=q�����2����_����_�|���8��!�X���]�~�t�?y�Q�����>^ԙ�_xr���������~����tm����t3|{����z�9�?ϝ�������������=?u����tZ���-�?_}A�G݊��������g<)���3�ޔ�(�G���#��g����w��t���yK@��a�ˠY�x��xn�	�3��M����ɲ����mz:�E_���_lX��w�����/~���?~�/����?��������|�_rx潇:z�6���&X��l|j\�)�OA:<�>]%�?���PK   L��S1t&�  ב  /   images/3a57aa21-29d3-4406-b48e-ea0158aa2049.pngԻeP�A�6��kp	��5��C����\K 8��,܂����Y�<���<U�����,����3=-W_��~Q��@A$@  (R�b�  �%<,�)�;�	�������'T� �H�	��?\r�V�z<�Yj�
�3��J!��l"��ʶL}!gE���l�����,_�!�EU�u\tT�|0]��p���g��נ�K����c���;-]ü7�3O�G����`j�G{��8u�rc>a�i]gbg�4��������L��}�97c��L=��`�=V�s?|f��<�L�8��"u�u��2�9����Y��V�c�s|�+S�s�뾒�OĖ������C[�C{�4Gx8�0N�ArزLbN�pK����e߆�6�~����¶_K��a���^]S��0�1i���CLi��E�!�[n�q�P\�bc"�X�cS��ԋKS���z{��G��J��^GC��OV�݌��u����֋M%���k鈿P�H��[�}�`o�p��o�M����Đ���F�ĳ�U��~���U3�-!w�M��!W�ȷ����6�3����ψԙ�5�A�����;DV��*��EE�����R���+h�ñ�Ԟ�O�.�y�oDQLH>"�D��SC�d�� �<o#���� ���t����MA�+2������JshBm���RB��À8�}��U��� .*�C~s2V�U���?��y����C�#:)� �q�� zfh�(62��po߽k�~iD���sG|���;<(�w��r�{ qoP2��މ0��(�¾wm��YO�T2�9��3��Ä��g:�����<��1�1�+v�p�m!έZD(��$� ��~&x�|��y�p���OI��=�_#���U���'{w�Q�A��ȗ2��6K��G�J6�J����ؐ��:u��]�e��2�^��R۲�L@���
�j�����G�V03���j�_�F �B\]��aD�m7��U���}Qw�"��x��s�M7|32�ù@y\��h.׼������'Eg;J�ꞣ�u�,�sy_(Z��w��\��Uoh�w�Z�u�!%�NU@mq������)��y��Î}-*�O�:��J�q��wy��Ah�!�3d����r��g���MƑ��pW|j�1&���3���	iٜqsާ��Ո�WCd�Gs�p�,��&y�c�pf8���H��[8�+�������4�]�{_fP,)A��[���;�ң����\p�W'QͶ� 1�5�����ȹ���l��`���%-m����U�Z�p��ДQ1f���ـ�vVCeu�Q5]������ҷ�� ��'�.��|y��ӑ���7��'0���p���vރD1�o7Mĸ;or��ռZ"*�hƋS�����������$�l}cA-�F�ٞ�/qz����r����>.�b����:�`3�O���I@cH���A��d�����{�Ñ���|�� t}	��Z\�6^��5v[�-�ͷaD���m-�-��z�����G��[h"A��z�������]�H�I;�U��ӥC��@�;���pA~���5� ��`�R�Bri*ZG���#�:�?��.���e� �G���|������ �����Z88����-���{���LM�LA�q�`2�������9-H�nG��^�tu3^�~�>c��-JP69���洦]��X�����.ar{�(�p�g��E���z�=ӧ�iY��������h/��t�͛�%VaLj߇x�ڞ/�n�D^-Z�m�f8q��ܫ����0��9�4���	f1���3m�o��(Yp�gc^F�-M��T��^�o�o52_7p=�v�1�f*�J�v�6s��yJݽy��V׶"i�j$
F����V#�y<l� #$�C�K}p�v�ٸ�ͥ�m>�?د����:�X0h�R-o��F7���G����(�4����ig��gq���FNA4Ƨ���KZ.����[�Ō�����#�֎Tl����b��c����/��!S��W�ޗg<�6�����[W�V�,y���=�\'@��)/W8�\;�A4%E-�!+��J��u�w�f��@�����O���N�g�H��W�ȅ��/��eův�[����:����Gl���.A���m�nύ�i�$l��^�r�XNU��X"�l��o�*�Z?�5 F��|C ����ђ��C<iI�\�m1I5�Fw���i�p,5C�6�Rc�+�� ;E%]�˧'}?�$b��@5C��7@
���'Zw�X���̞@��P6����>z&�"g�ӑ6��I�N���2�{l50R��Է�G�5VW2Ǫ��AW�3�tp>~m�+���W��r\-����	Q3�h�mU��/��tڕ�y̙���!�e��l[��ɮƧ�%*m��:�����ʴ�!����X=�RHB�Ɩ�?��	��젮v����Hk>�"���,�A7�~e�v�Nbka�2��Ym.!i,�쌍8�u_U�i�F��F02Y��֣���v��WC)��$"��XگPq�j������ӌ��VԀ���3�9�w��]1����Cmvɴ��P����S��pJ�HX��{�d�U�(��QݜB���I �7^�t}I}���@8G�}.R}����EI4\�Mw��cGc��'y�Y2ţ:Yy#�^��
�|_�$]nP��aJ��U�=Û�t8""h�}{������&�]���
���%^���䙆��8��Ee^���@���Ŝr��.�� �>�'�\&��Q����}�e�Ҙ��sMu�I��aN�~F�i�~e�U+K?���4[|�s8a qW���!Ƣ.�b$�j򢴼"ks,Ѵřoù\�.Wqb�6��w�*G��sC�؎�fhI�����]�ԻA?����������~V"~L]�F
��?�ʆkko�gq�ߟ�8ѱ\��EJ���a+�s@ҰQYD����PbG%ⅉ���_Z���y���$R��	Ë���1��}eG��г.��!�u�ǎ�%���P�c]��y���[���M(:jw]��	QAs�<���j�(<������@�ʛ{�xў+eۺ�	yڈ�:'����j������5�Y�7$jS2i�x5������O�N��^�,)��f�Y��A�IK^_�r�6>��SԎ���L.\)��N�f�ʂ���[#͍������j���W4�V(^�����������X���tn�rKo�xfZ���ԕ�V3諟�: �{��+�\k�J�J�vZ��D=S��ո����9���14���t�^~���%��0l�����$���m{e2�0-V��G�Mi�WQ��2��g���2�q��g�M�,9����4+T���q8��j��:%�vCi�[or�UaU�9���{��N�&�]�W��~W\^�\<���t�>�o�xI������M�$du\$�4�����L�3p��%��Dk�I��R0���î4u;�@Mc���X|����V��OY#5ET�F�6��9JtꖣH�@m�!چ�J�ݍ���҉�l�J�409�|��#�c�Q	���n~�ys��8�~~��F�~��:M&y�"iT��UB�QЀ��eNS&���5H�,-�t����a�����۱��ě-))>Ӹ��R�����W�2+��2^��8o�%�~ʍFPkvUdoU���A��\����C�������x�L&���w~R{�i�����w��^cN�]i_��Po����Ԍw1���R|&Z�R,W����|E�~��7j���<խ 5�Rb�0�.K��@Y���J�Y���q�'��eRc��#U��-���<�-;d["nE��� ��	�d�4�[WJ	V,1��RZ��"�g�z��Q�s�NF��O��\��]İ����[y��C�<�]#SH[<#C�+�e�7=�ӕ	=Ѥ�Bg�d�S�3�ru>���ݕ���/�^��<�H<AI)�A�n�4H���+�e9�Xc�:�w��!c4���l�h4B	`��j 8oZ8l;T<`�p��(sME��,;ӐsO�L@˃1�M��\N�q�;]�g��V��5")��F KE���=wQ��
ov���fsu9\
�;�۲T5ޚ�W@��cgZ�{^&И`J�H�S��xw�\�⳯C��~J)�QN0�p���G}�����^��'�s����e/h���ƙ���"�Q*�T��6Kӥ�i�2��#�i��f΢{Mu�]ks�Q~&��>�O�u�h^�����+eiO��k&[��Y��.|��0�f�D�V���}`|F�ȒN���U��9��gXSዧ�����������:��O�L`k���Vg��B[ԣk]e6_��jNsinbWY�O"��t�?�}����>�җ�A�yX����x�ԓ�0��7W(�	���=�c��me)i�y}����MΒ����:���ѽ�Y*�W��<LW_~��FGY���e)W�Vd�>���e=�㬱�"����n��VIK!����3Ej���D�1f��T
"�g�k�{tW8��>����\+[;c�����췬1�Y�/����bT6��k�8���e��YȾG��5f�'����c� ���)ޓ�r��7�_�d?5���t�;�B���dI���N�2��S������ת���]f�L?|�ܭA�����N��7�V�������q	o6N�>��ϧ�T�Y����c�Fs����K`*oЕǃf���e[��lYN���y�3\�.>�U4B*:��`Oٝ�u1�խ�����E���f��/��x��Rg�� r�j���՗����k@�.�!
9�9���r���F����;�[���&��RuJ����-W"sU>��S����w��j�����:���6�&-�p�Hl�mϿ�zR�,hd���4���1cq��~�.
����v)h�ݟ��ak�n����}�q�cw��)v�.E%.��s�į�O���8sUh_��S���♊މڞ�����t�\���rHgҸ��@��rE��!���{�J��\���t���?�I���q"zH�1�G�\}l��z�Jet����������B�N��	V�g��
�HR�`Q%&����}�<��/��#�7j��k��:r��O�o[��Ev��ܽP���*�O�NM9FLX�fA(a�
�s%�ʚj�BQb|<�|,�\!��<��U���gϥ�}���
�`Đ�wA�6!�*���wߙ�=]k��m{P��\��-�46m*G���M��9�� �]4]�x��[��>�/�u��N����9B��y�4m���ٽ���Ul����P��$2� {Ѭ~�@�lͱ���r��Jכ�3�t��^����e�Yߐ�չ;e��C旍����էo��iz����\��_kx�{��W��ߑ ^��S��`�O�a��Żg�_��0�D��S�;،'�Q�;a��C�87�WW���f��چ��Պ&���F���t�O����5�-�WL8��b9n��g�3���P(��Y��&�Yw��*t>���}g��W�����_&���X3	�(��i\����w�p� pS �֥��k��_�	2@'q�x�I9��Q�[)G����Df��VK�c#�
�g�"n�U�S�����דp� 4@�g%M]���@�=j�p�gdGEf)=����t�&��"��q�)6�w� �/扩��{�ݎ��������}J��
�4:Վğ�a6,��Q���u)��d��/��=D������s�0 �}�QTVQ�r�'i��Q�z�\Z��XW^?[TqM ����m(�<s`6&#��N�?9
)�S|�oc�/�X,�B��"}��*�ٴSR�f>6�&v�P29�څ-�|A����2%������ �d���<BZ���=~����`��3��v� U���&v�Žx>�5맮�Z��g�t)�~��������T�Wt ������/躌�b���A;���ߩŕ`9�XD)�Ϝ+���qX��x�\�h��.�A��~�����g�}��{�y�T!�{J���(�i�dc��3��>��O}�t�Zݱ�IJ�SF`	ylm���88�+~aQ|gh��'�6Y6�d _���O��@��l�{��nJ<���+Zo����|����{E�1
5�a�`�[�5�p��h	v�}�Y�A4�-�)T�y��o�TI4d�c�6D��<�2��J�II!�ݟ
A&�S2S�]I|0�A���B�l�ص����d8�4���O'��y1�� |�=_�ӓn�
K�ś���y�8^����ݛ����"ȱ�S2w�$a��fΌRqo��:1�~�f��r�	Ѩ���ޭ1�����'$IO2�7�BZ�};C��O�L�Ǔ�xߒW
�|<���cT�~D���p1�߳�H{����!v����ɘ�Ln����C:{E����r�W$i�>�����H[48�3]�����@�[��Ă{IB�U���+1���,w���-c�妠z���Lp�+eJ��!���E���E�^Տ$"Ὃ�*�׊Ӡ�DD?�|iQd�/��4;����JW-��Y��v�H�/��n�XX���3V��r�OLyw�0X��z[�����qU���p!�As��W�iIt 7���N�7D��s��8�z���Ԇ7�w$l͵�|��<�k�&�"w;
�[T*�T��A_�t����d��-��)��!{�
Jce����lX�A�<���bse/,��ҪX�x��ڔ�����
ɢ�=����(%���7�>= �YE�ҫ#�Cz׺������^��Y�Zr��S�@���T`0)��
��;���?V���iA^���y��m��/��p?�*�TK2��Qc�*��!�dh;�IEXt"��w���
�߅ɔ�|�N8G;@f�E�?)W-���K���$#���3~�x�#"�k](����h������=OT?a��]��m{��U����9veh����Y�[Y/7A���%ˍ��|}q�b_���@WM.�z��$h��(LLy|��}�Q�����"U#�
S���G��b��E�[33�\��� �>���I�:���[6�G�]����¤�>��Ϫ�]������i�%�'%p��7���9tF��+���o�?+2�ۗx��g��B�&h;�S h�Ͻ6y�TT��`R��M��Y�0��iѿy���&�(hM"t���Ù�S��d^7ՂA=���&l=q�~�O��T��x�d���=B��ǉ����w'�HƋ�[���oJΦ:*��~5L�%��r})B��&_�!l�+�.�.&\x�p��}T��3�J�q2<w|�Nn�;�f�n�V�`Z�E������u������f�r�HD��g�F#%���$�v+u�X?���_�K�'����8�&�qM�V\웩V���K4
ˇů����3����8iN^g<C�U�S&^j-c]:���R>y��?T�*`p����A�Km���"�UܺP��}}��P��u�f���ڛ����ү�o�@	�0��f�9�(̹'�Et���0�x���6u�0fl4aL.ѼC ,@�2)�s���'��mz��-��sU�oL��Pg\ZP�G�p��#�O�n�V�ޟ���tX;�~NTگ�/\_x��I+��]�}�خ�E��9��t�{�&|�Z�m�{�eW��*�}i{;�Mh��0�q�?��p��5{�K���&����4h��9�Oe} ��M�X�����/�C�����9?�����XȤ�)G�Y��E�^�s����,�n����H ��B23��	�h��.z?��s��C�cpa��q�yf?�w?8�t�`��mF�!� p�#Y�#㿔L� �^�5��D�)V�����+�rO 4��9oH5*B�ܴ8KS}L�W���yP�qjY�q�'�}�\�Y���v�A�N��ajPu��P�t��)R���߅��k���_©:��B`Tpޞpz�����$2�	�/L�6�4[��5�
\3�{`���V�uMp7��$���i'}��V�Y��|D�׹�>mŉ��|�xʚv�k�:��Sp�,z�^�"�T�Sy�=����~Q��床���o
�32N��q�V����._�j���⻈�j���%�d�%B,�ʬ���JF{��F˅}�@��mx���~�Zl��۟�I�Nwd��3"z����iIV+Vj�Ϧ}����u}~����T_G���&�2ҹ��1���y��h�ZT���h���%34G�i�o��f �<��?��Рxyg0t�A��5o[M˼߫�#����L	�A�� �py,�(_��Ɩ{{���<�~jFi�6Ɂ��(j�	2�d)����f�.hغ��W�(%�k�(,�/��ېXX0j�u. f�V������@<�5������,�wm��q�g���]w�E��u-�_u�׶�SG<d�z�nnRC�ߑ��+\Q��"�t��Z<֝��ZN@�KC�#�O-[f�=WJ��Eo�������;�9�F����#h�b�-s�Έm`ɳ�DF�ĮY�D���\�(=�_�uq�oN㽒�' ��e���^eegGݰ��w�Vfk����[-��x�V�l�0�E����gƋ��Z�IN�G����V�ۤ9Å�*�u�K�)�[�y���K��[��Ԋ���2�i��e���k+���� �����(�#Q��V��~Tnq�d��(Y{Bu�t�|����N��B�M,e��;�Z���1k�v�vؐf�9�d��\�}���e�Fbl$R7$�c�@�"WB�<<3��F��MDܬB�#~9�(2�Lp2G*�M^��*�9*���~���O@��5*̅��I�
�S����N�#���g_�m�F�|-n4��<|�p�_�RՓ��񊷰�fs��o�F�p6Sl�VX\N
ٻ�4�{.����"MW$��n��:�p�",(k=C��MQ�j�
Ց��y�jF��p��M]�W�K�+������|ox�t?Fع
���ٞ�v�i��I�,���tr^{6�a/T9C��U?J2J�躐�Y�N�43���C>Q����]��;IQ��i�)6W-%�4�|�hE~y�E��Y@����	��Eϭ����7�#�ͷ���x��X?v�
�]͒pEP%ց�~g�6�6��g��Q#D���N��C���3ƽ1ݕF]�V��̭�@�V�g�����jyA��� Q5�Fc>��`"�+4���DY]��:��a�����Y�����������L��� S�⠐�g�)~��+(���h�M2
�c�ƒ�64� ~E���	�>Y�	 ͓���iWI�^�ԍ(͘��m2U7��x��i`�t2���<*χ�P�>kŪE{O�e$�)A�l����0N|�����j����/e]��`5)Fត/d-*�N�_�g�Mrc�U�Q67��
�^�K�E�<�v-�bŜ�r�G�M�k-IŎ�Ǧq��Kώ�udX�5�6ނSѯ��i���yכ�ػ]�Y# �!�����hnt��*,�1�U4>�9�������*Ֆ�C��{�x4x�D������Q|GL5w�����%�$D�O̳UC5hvV�
���!��k[��*�4Q()UjSx�2�|��:X�QO�O/��z�@gX���㧞���VD��e���Q2>���Y������S��0m+|#����8�C�<^ Ē���o3�KvqfG��R@jKw��"0rԈ�$O�ҁ��a����8��Ml��6�9�`�������	#0V`޲l�ڭ)����^�^�D�٧��g?��$�7�B���'�k���Y�W��:��vb��(Q+'E;�r��K�v�6� m?Qd��-��U�εQ��UQ��Q�a�z|J����I�d���i�Δۂ(�f�wQ��1\%��h�`ooE�P}��v���'f,󈨉O��eb�㰹%�%b�S��sd]אfx���D`9�D6����!�,&�E�x+;���"��z��_�vY����0�5��/˸qUt���g=?i0Pw�	�<���ފ#�r{~J���������7�,��<�)���t�;��P㔕�����+��Lż��3���]<k�'w�����񮪍�3�̅�ÌH���Z�W��	���c]L�˼�;��0���Բ
��!^����.ƋuS�����2����s�t�����!�zO�|6�E31w8c��`���ˋh����-�~ٓ�^�y���W�� 	��q͉�����\g�u��g�<���J��4��s~�OPI���%���a��>|�E��[Kn�J,��͌�m�w>��G�^��Pb�3ۧ1A���J�!~�A|)�l���[�Ȯ;����n�����I�#�oG�߈�P�S���r�.�@��a>+�~k�0-RY��e/ۇ��������	0��p�`�����ם=�͚ǚ����}�@������n�(Ԓt}��*ǿT�:�;j��9JG����v�ԁ��]����n�S��[�n�?����f�RO��e��߄�<^ʿk����si�� {���L���o;v�J�Rj����m*�5]F�A��j��������@h�@B��2S�{�1(�>�9���W�:��^{�q�IK��w��	�8c�^5G��e��h�t᜼FA��s��s�敖i��▐=�@�����R��=��]�1_����pC�R����r�d9Y�d�vډ�~֍�=�����\s6��d�[�}�J�d."����:��Z��e
�tΘ��Jʪ֟��=!)��HO����j��\hL��Vn<�&d��=E2PH�@al{�.ni��'����w� ں�q|��'dtC�N����s�����ߋ�LFw��'��������݇�������Al� {��ۥ�`� /��$[������dq�=v���䅙%��y� x@�<�+��2a�gk����X�|�q��� �g���a����*(Md�����9�ӻ2�����gD�q8s���T=���h�D	I�p�x�עY��,^s��H�nV[��)��'X?T�й��pcOS��DUu�~��s�%�f��(��"d����%���]�q>c-�%�[6��q%(���m��:
��\4V�:R�3.h(V�[1m���_���׉�RxL�8���<9�"e�T)3��*�L������{�^p�=��9�Knz�����A:7�^B��@�0%�hѕ�\�Y��#����ȕ3�=�w��W�mp����LX�Z[o,�#��=j*�!���Fw��������A�jV�.^�o���� �fn���b���@��e�Ӗ��ˢ����8aQ��:�<�=��4%18���3�;i�}g�6Fk�# ���L��S����T��˭�a>D���-�����FGa{,J��s&=`b�Q/�:e���	��rԘ������a���g������`�ͬ��l�� ���s�2|ʺ���}���2E���m�^J��I�im���I��,�+�_�Ҩ����٣e��]Nr��%��6;�H�2O&@�j�Wۦa���%���D��~#�m��)u��+�G���̈́��xy-����ȥ����@e�9=�k,~�M}����D�v(�����-1�o����6�Z<�M|���!��`u���9�͙'�ԝ�ݶ��П\
���ᩰ���!�^�n���bT��|k�jQ]O�m���lpp�l�<�"�<��9�I��G�	KH�ի�QKֽzKǈn�WMm;O(�'c��� I1��>��(�9�9tq���$��Wrqqǰ�L���c{�#��a��sFMM�]DX]��X��;�wCX�fh�$X��*pw�Sr�6�g<��,Z�M�58��3�T����}8�~5Vj��c��i�S/��ut����C���d��i�}Eo��{�f)sx���5��¼3�T�ҷ?����h�xH�1�-���K��F#��Nm�� ������P11ƶ�+;�l_r��hBP	�]�]�"���$z�-��IƮ��߰{�aj,S�P
�D�����F��r��:�A7�4G4&���4��h���{{Rٍʂ�õ*6C�M����e��� 5w�ڼi�w� k����77+~�9�V��_bc+��s��D����t	�!��?��t�T �"b�w;g��'2�>��'���J�]����M�+��0���Z�5����&})>�f�K�O˄��P�h�#����l��h]fM)7Љ�i��s�u���<�:2�uH��Q�r�I�jcI��a
&�vG�^e*��^��������Ψ�憆�����(BNy�qz9_�`��RL�l��R��c�6kF|��0^�)���cV���.
Ρ��!�����ӷ�	�/1u���v��p]a.i���� Cԣ�.Y��F+8����nF��� �d�oi�`��dH`i���������N���G����E;�67�m�m��b[�b)o�|}#�p�����@\�)S[���T�P:m��+1]�����O��x���*ט����4T&V� �!N)�J����j&��/<��IG����Q~&�G�%��Y�Ƭ�g��Ŵ �f,���s�������4��mOy�d\����܏^��,�L�z.�'���Y��rV�;�`�]��	��V+��:���>{���/�����:C`h�kFt��ßklK>���Lnxg�	&�\�i�T� ��K�@�Y\ڔp�:�q��b�z���|F�K�Uw��j괦t����WngR,	ah6-�_r�=�!nW�_�G�S�%��������鐺{%�H՟�k�~NB
᳀� ����{{��ʆ��J2'L�����Af�:p�>�Z��,n��.,���`_y�6C��+��*��㒐����ZL�w�ю��]"0i�����b��p *�=.Z�V��?UWO#ۿM���zh�Г䯬e��I�fc��1�?p���s���T�?6#�9*@��E('�a%/4�Z������v	S��_�x9�c�G�_�૩֙.zS�� u}�ũ�fહ������7<!�ZC^�-,� �Vu��h1��kW���0d&�-��ʦ��*C�y�a4���u�B9Y�K�� (
8�M�q���2������X�	P\j.�A��tܚS?�sQ0$�^x����T�>�[�������B�]Uհ�T�.}�bZ[�B�E��/��z��W�L�i_�s�O�oo0�"a Q��v��Hh�^TCI�����,�c �.�caO�ۤ�����]v«Á��Q/fO5`�C�X:�9F��酓����;�! ��6���B�g��Œ�ү��J>=�j�7G�w�v��{xOg��,�P�e���/#�ߘ1)S:U�?�)���~��� �	e��Ƶ�(iʄY�tqj4[N6�(&��z�� AR=�sMv�x�Aw��f���[�7��� ��4ѕ���gM{w���_�!��-/<��?���t�Li�p�uw<��F�vV�,��O��8V�⽷1FŅF8�0K�Ma���X��hp�.sw^˥rŅ�/wU�:tu���;����@��$�"��g���r�|��=<�l9��C'�ů�0Pe�I�BX$�����Ol�*~�����2d�| ����|TY�6���./�R?��� ���{�������>��4K�v�2��!��w���ͪŮ]���4k�����r?������5� S� �W~�����iO��L@+���O���V<��fb,��3^�Ͱ��UĪG�|ig�����+���yc��.xg�=����ՠ}Ԇ*0�j�M}P7��2u�������/��vF$�bEGW��=�Y�%3ڢ,;[�7��>:7�=ӏ	�K��بd���IH��ʭK�R�*0z�z�y��b8��C�_��$���l���.�A~��M�� gE�	� *df�[`G�ٻ�#�#�(���_��+͡3�6]�K{����f�(���b޼};�n��g?�Z��1Gp���'��yh���qc�Pc!�2;����	CL��î�����ڈ����V�l���ۘa��B���Z	������Nw����� ���˺�c[�\7i;�a���F�^�-k���k�#������`��fz��]9�7��m����[�����&�G�(�%�5d] h18Bs�0t~��3u�^�N�Q<(ð�p���L��s`�9S��c�Ɉ�v����+O�}�fj���fͭ�xz�&rB���]_Q���5r)n㫧�@Y�ꥸN.3�qYo�)�χ�?h)��z�L0��/��������qu��4�O������6�~xc_��*i,��1Y��ZM[�
6_�u;��W�ŚM>�U�K�=�����Gێ�u���o�#����\���g��b�>Z���&Z=a�6'�3������M��ڤ���I�M�
�s3��M���g�����LT�v��v�����9�ur��9�{��I�^L'�t����wn˭|�!�9�y{������o%�_(��>g�;k�+��� !�H�a_2`Bf�y�s9\�_Z�{y]\�\�J4��kDN��� O�sd���W��G2ds�X�4� �a�C!�]W�%H������*/{�'�Rڜz����ءzW�"�G�D�C?�+q ����G������~���W���T��!����� a��Z��TƗ�Ǉ����T���=0�����0g]�-P���+�.+���T�j��?c����~�=�����Bu�^yX_��"�w|��0!�_%���]g��5h�w� )/�����gŭ��3���o������:r��p�ZB�0�ɨ"�Է�=fv$@����_u�Y�j�^�m��n��vc��qL�>F�-wbZ��� c?� 	-vUx���^;}�X%QJ��9�^+١��ܤ��s�l�b2�D�h����֜�%��%T����Y'��U�F*��+u(#-��
�\��q9r%n��*�>fj��Z�b�ײ)&*��@\�-ŴrsԕQ�*(�0��e�C* )2Vdb6Mj����6י��yM�\�B$w�ZVR6&Bql.��7s�j���E�����}��Z�?�ū[�'M��/�5n��|o��q�o���q���j�<�7on���o��z�#X9@_�P��.�Q�F�� J�v��T��K�qӷ�ֺ��T4�R�Z��n���I5E�u�yu��݃1m��6u+��f����3���׆@��T�-/��rM�L��$d���eM���VE�֨֯���}Y5����#.9rք��h��0��R�,d>h�Իa�m[ϖ.&��5tJ�Uc��"$+��Y��0p����p�ɋ;�R��L(MD�M7U7�B�L��&�C�5�Zd�|d��%N�s	�jq75�g�0��.�
������I<FDXw ��w�I��M����w�_�Ƹ�)��ۚ}�Z�����M �5 ��#Y��@Gn0�õU��8i��C������}�\�"���ξNj���q\D�o�o���S��¹����w��iP6��׹�zs!�%���c�q������*s�����Ƣ�1��9���T���3�]�ll�W� }�HIM������#�ov�n��1S A���=��\#���b��XKf �G�y�	��������#B���A��<6��;��M�B�G����E��Z�_�m���G�+��f�[s��[!A{�h��4���o�9����uE%���@HM:�_��]f5!�bz���o�JK�� ��G�Ʒ��LIII!KK1%1�}��q51X����r@Nn.��?G�HII1}��3�WSS�f�A���G��fٍ�c�z�ӆqY�k%+��oG\�����)9s�c��k���А�������w*~�OT��(*������:*''��^���������7Vtqjjj���,7����}���ƞ���4*��ʁ[1


*ZZQ]]"�݃�����`����웗0/�7������Hl�+���ߞB�L�R��*��֙�GiRd�/10��+.,,�
��`IUU,@9j�k3���ߔPB2�H� $$<fq��-������a��� 			�\�H�;4 8��J����a#�*b��_Ц"$�CL|III	G}�Go-ob/xt'�-<�J�ta�l�eI�7	?�͂���oWOZ��Ÿeϵj�թ�/��߹��#�>�/~<���1�>>��G�����'�\��5��5��ݴ9ɫ]y%bJ�1M�O�����y��>A"3!�%Jřr'k!�w��kQD�BAϑ��ǽ���h�8��{3�QE��e�%%e�9�x�8��{]F�kS���J&������gs��7  Pd�@?�y�`��49��Ŀ���i_���,������qC���ob�8�Y�a����
#�T\,�7St�#7� �>��7��Wׅ�����7I ?�̿��P�q����0c#�e%�N <�K�H�,�:��xU�u�U�W�2��f��kA�g�������6a�7��ndHct֚;T���}QЙ��[*�v�������o&"�ǎ��Q.1�n6j̳=��f�G�c7��\������7�y���Pn��c��l�3VFG����3�������`������H�W��U�Hｾ��� ��H�J �" ]J��� $�Ox����~8_�g������U��7�z2�q>x���ݭ8C�h ��*aP�u<�,�zTI�ܛ��jMF�
%²��V��l���͢����9��8�|�.[�%��B�]y�~Ŋ��oؐN�©(d��K&��ڭUq���=��fo&bt@_?���e���y'ܤ�������̐\�%%iv�	�i}_y�����9؁�[r'�����g�#}I��{摐�V��BS��� �.�I�;���	'x_���u�6Y&���f��#bW�'-α��B�o��vɕ���/+l���n��OP���b��K�>I�ߙiJ��!`=�/�a��
���{G`����r�������'���(�]T���d�����b�A�.Ny���>k(	4�eF���ߜb�ٙ�Ӟ��u��0p�\]I���M)�~���:%%�K��S2p�0��|4���+%�WohZDJu��꩓5T�������ERb>�4�F{�Q᜸�g��
�܉�9mq��"��D����$RA~�� 0�&j:�f�a��Z��_8I35���Yur�$e8��[���K�����C�s�Y��Z&Y�F|A�`Ap��T���F���9fo� mW���R��O�����ޚ�&:s�v��'O�?f���[��X��_�p˦�G��ܲ��8��KE.\uv*���N1Ix�`��͙('��'z
ހ�&])a�꒮��Cz'�c��i�}�X�y|��%�(*�o}�0���0��*�����'L)� w�S����c9b��B H6WQ�OаZ���������VD)�'�֎]�ۜ쉭e�zvlj�5B��bvn����a>O/�n0-B�M�1��Kzs:���tl
�o��J�z���էJ_>iw�!�X
`�(una� brM��^�-n3�!�%����t��������pv;���*T��ARd����2W��`�r(ת�;�#{d_� ��g�F�c}��������g�#-?�����ޖ�I���]C�r���S�X�i�.�K� ���#K]Ë�tT�����6�fP�Vm��RK�<�?Ġ�64T����C>�9�U�kB=������N��Z���A$J�w:U"P�H��e�{�V�"��D�?(�5
�v#0����ֻc&B5���B"X�XZ���-�J���\����P�Z��yƮ�C�)���NV	���i]߂R��F�}���a��!:ҏ�5��R��4��p��z��fJ@�I�0���fm��1G�K�"c�!�4��o�v��,�{B���|�Ht�rZ�W��G��U��|P����f��|�Q �6�V���C9��z>���Loݲ7���	FD�ʬ*L2p��8�_���k��x7>E!���~�mM@�kf/Y�3�»m9���*l-TЛ�����HAk���.Y���DQr��dU�`��6H�κ��3�	f9���ĺYC0�����e�B��ѦT�o~*1��=}7kAw�a]k'�e��
�ZKސ��>�{o�����Vc�~L�`�PO�i�nI>���/a�|Lɫ�:�%U��2��,���v<6��eq����Cdݧ�4]�.�*�T���.w�W;P�ޫ����'D����Ϛ���;\��hے!�����g<�5f���<Qt�� ���Հ�>u�MuP�Y�8�%=~l�ũ�^_��Gp ��?- :X�-B���+���8pH��$JXDW�����ӿ�L�|���"_�]���:r�N�k����_8x�}���Ν��<��-q��-}�~r �Θ���v�8�����9@��hհ
�OT��<�:t��]��:[��fR�����L���
N>Įd��a��[q;�Ji��wbσ�A�s�	��:�Pq��Y�iSa�H߃��te���X/��#�iԜ�O���:r+�
z�C���N/Kq �o;d���#�KX�Aaե�遪�{Y	[?��;���uL���mM��
ڐL{ �M$� ��N�����g����`H�J����;Ï�k�ָ[ິ����P+X]W%W�v��Wy��}BZy���]��R��'aT겞B�t�֊��t<b��ޮM;ٲ1�CGQo|���2T��B��һ�}����f8�
�-��+b6D< ����*op���� &=�zHF�&�\Q�R��\nJ�,s}:\ѝU�6T��kh�=���A��N�h"�p��I-H)XI+.ш\�"ơ4����:ʓ?+Ry�o���,�D�p�?����.N4Ȓ�'��OQ�i�A�BG�������!���߶P:�Q?YZ�\�,���͕���
�a�G�n[�n[K���:-�#$�' ̗����I�%��zܻݶ�3� �/`%~�T�B_��%Pη��=^q����Սv�K���0�=sl�W|J�</�'nӪFu�g���r[�ǈ:�D��,>a��p�;�:�;�������u�PWXp��:ڲZ�1Z���MغZ��fXt����}X�{Oٮ�J����P��Ӱ9́�qzr{j���e��J��߃�����b����.iC�N�V��r�X�&Ĕ���������;`��nL_d-w~���34��l������6_���-���X)�Ț'����_��W[�1�N�õ�.1��G���'.��%���,j�� #����5T*��a |���O:E|�,��B~�m�,�������Q��4e$s%��������z�4�`s�E98����o|�y�wh�%�?K�e5���
��GgO�8�z;��64��Uύ�m�~�Y��;f0���7�p�L�$p1���lw,<�~��%:M����7M�;���ǰ��-E�]�a���cKhߛ��l<D��?��~���``���g��}+�$&1%�Z���e&���8ܑ��CF7��q��v��A�`�L¡/e�U������ZL�0Q���R���z��vl�����S��{��)�I6-��!��I6�nO�����يYZb-I2�-��̃�B��_<�P���!�\$�#�ny��LN;������r�d�P���%�.�Fu)��c)k���E��=Z�Jsw��>����N�m�`M���D��:ÂGd�Ӎ�}�N�":���L��v�9u�}��N�{�;���^��r�F��#B�zR�7B���_�8�'*{�����1ֻ�i�%%eb���$��7�)���Z@T��z7�;U\k��f����4��@��ғ]^����+�TX��1%���E�aXE�q��4[_�]�~�Rk�8<Pș9x� z��ы���5A�둈a# ���6����h`�]Ʋ1:��uw���L�ɐ���9}����0F�ro�M�Hd��.��c�%k�r���3� Wb"dn-� ��?�Sƍ�,h$K[z�A�0�>��#J��¶��k�㺌v�n������}/w� &�3?Mo�˽�AG�V����C*=n�c���M�!�T�����A9�m�2����]�I����3-�^��Io��gn��,��O�J��UP)���*�5����$u=�P,U&��8t6�i+W��+K�\Pbm�k�gai<�8t!��&�����)�o�h��QO�bm ��Ɓ�c��48�G�3��8lo,��&x�f�f�9��I�[��Ff��b��9�U��F�.<�p��dd`Y�S�UP���5�������B)�tx_����[2��9�4�kLH�?���=�iL�d�ɖ�$T�INЃ#҇I��+���Hr؁��J)����>ߍ��~>���29B'���:u�p��B\�Z���)���I�mP��)n-~�j�b�/��olF���L��j�9�a%�`�
��l�����^�F��=��ʶ%�-n��P��&�}��l�;���:�sӒ%"���deK�57s��a��3^@}�u1�6k��K�{l�z�A�*=7�t��֌Y�kXt���ts�@�/����1�u3��g@.�P{8��ꮂ�K����m֦���Ǥ���0N9#3�"��-bz�?� �3p����{���؄�ǃ���|�ä1�� Ec���ݚ��t`P�{`���ظ0���d�����)�T��%�*(3��.��e�� �F�Φ6Ibun=�(�2{圽]����_�l�? ���<U4o�O���� X��$n���?�c�Г.�ĸ�"�B��>��x�T԰�g�"��+;�]$Q��Hi�.�X�$6�� y�$��|8N���j Q�[�^�`���E�Or���L��&N������[v�|r��`����&��)ByK62te�F�z��8ׄf)��f� �Ja�p��U��E�9~�`�1z���%>g�.��hY�-�q��`�����jT�I$������3R� SX�`G��=B��In����j�:�����"�>ɍ��g���x���)'��a�'�R'��t&����[c�! ���Ty*��jZ�H	$#�K��co��Ks�I���vg�x�*̹��/����'�	ғ��ݾ�{�M��@��p��������ey댸��c�-��Y�P�^���VoX�9���0�
��1X�%'�09�#��ʹgWVu�	��X����t�O6��(������ig�q���� �kB>s9|\k�U��b���]�Ȓ��O �	�Zw�
ᩂt�;�b�<��Ź��OYt����y5d�pL�M��}37�$��������i�m��d��|t6��9����Ҵ�NHt���lv�Ga;�.{n�}��� �/�F�]�S�Eׅ0���W#6,�\Y��:����ӁuB�m?���SM�d\��X��.�2��Z3I�}�ۨ�I�m{�a��W3S��!��u��!#�qq-�~��3q����]j�r���Ϫ��!N_��C���Z�]'$�,�K��E��H��rB,�,��.�K�Xќ3Z��{��WE_;���n|�MX���7+ߏX�B�hA��:F�)��X-��w��SQ̥�����p����O=~a��{m2��ڵ�b�-��🤫��G�dEw�����n�Gvj���n�B���N�@&���/�T`u�E�ڳ�(��3}��̜GE�y��p���	#�*���U�#�T�����r��5�G��=gjtN������}S+�p�KF`MLBH��,?ga�r�*�G�����8�1�\����P�XB��!�pu�����Ҽ���Α���ug�����H�K��\<��gwk4��pw~�7��&�F��b�;��wl=��L�a�"o��&SF�U�Ԧ�Z��^���te��ڜf]>]E�B�}6��s�O��H�a�,H���:H\�?�+ݨD��h���{5���_a���d���#y}���6�w��/�����Mu��	)&�k����i���s#�ֲ6�&��1A���B�Z�6Ʌ���#� 4����B�~�S.�.y`��N��ҩ�ob;��FP&�a�<ݟ�~�2N�[{���I�Ox�O,�^.i�;&����T�{'V��9*b��㻭�DR�f(��Ü�%% Wd��_~���v��ړv�f�\O�@\g]R��ZNkW�%�t6*�k�zt��w:RC �����J�L�r���O�[z�'7B�e��j.���	X��&Bc���v*喔�Ũ�z�o��^���7���e^?d���!�s"%��.A��BBc��ѹ����1�$z��%%I6�FU����ʑ�d�%��g}3k4�ٓ���z������p8��w�#��M�$澻�[]WF�Pe��lp��?����5��Pˣ�𩪀��j"|�G^��d�F���%z0kY	��T�����l�[��d?u]�WF��_AJ�O|�^0w�����޴�O� %�F��CC�߁Gx�0�����qY�J���/�	ZUu��b\,P�:�y
	/��O�>f�
W^�1��]��O��O\�l��LN�����huB�.x�Z�g�.��֬���s����}����q@�
xVTTp��o�K�I�ZF�38N��Q�|��7G�����Xy(nttT��ng�h��S��B[�%z���;��qz0����y1Iɜ�5��L��ht���<b}�����K��ZWt����(@��4O��XSccz��'��n��2W�M���+,�k�D���B_`�E9 ��xJg�|�~S}}}~�`�Z�9�����i�����̕��%Ҥ/����7���J #���w����7����h�[�����Lg�?y���6y�0$!�@O�FZqճ�5i���V�y9�n�Ss"�A/�v�	��-"=��car�!�k1���b�BZpء��U���փB	��]��RB���Ҁch}V��<�0��Y�Ϡ�(�l��",Bkj��5��9�2A�� �~K�Iɼ�����G_g���w�A+C��E�Ʀ��!Ѥ������(Eka�����I:F��V�7� d��p�jL����&"�l 8D�<���&T^���1l�V�|�ߙMI��,h�O����xVw6sŃg?H�>/�ao-�B$2����ɥ�!so���J�%.PиO�E�gء��턫��I|Hг���UѪ��r��}��+��G~��r+��i���p���,Xh�Q�t�>�h3gp$
�v��r&"��s�ŏQ@$� }n'nq/B�,��WC�fß\%���V���=���K�x�W��k ��=�C��Mԃ	�x�ҕ���>wR��G�O)-�d���@�4)	�PdL w@啎�Y�j�>��"��<H���*L/��~���U@;�r��(.ȹ�Q9�6�^�H��[KP7�W<p�}��x�P��)\!/@� �J���h�4=�J�T��##�M�����R��M�Ĺ�nL�Ž���o(mWW��~�79�H+�6�d�-�IkmR]��X�&Ş�w������g�m���<*�`xǦ��b�H��H+�ƚ>E`�(����e&(��Q*f;�?��n	j%�Tx6g��l�N8�ww֓�V����iL-ފ��=K(DS��2B�,���W$�X���|!I���'6sI�#�$�!��t��ZUX/0� f���m�Z��AaξK�X����� Y'm[���Y-��A���bWe���v�{|m|���gQ�c47 ��z�K�4�8։Å(���G$,1N����y�u���A#�t-��ѱ:�1�!��f�������4�?�5�ު�3�%��l����-��\�#�ex���l�a��GoeR�N�mzk�h��xi*����۲m޵�Hn;�� �����7�Z��z�^�JU��F�M�2�}V���hE]�:��-a�k�'���v��]���S������F�4�!����~nd>hUn�j��1v��WEnM��6�/d�SY�9�0|�硔j�Fta�n�L�W��
}Bi?�y��42�6b��F��WѦ[����/�pū�3En�nN i�]dծ�M|�"|�����!����('��9V�A�>ܖ�_�����F���u`�l��+�B������(|��9��Yڧ�}Jdm/����.pd|t3ARP�,�
�T���AE_����H��3�d��E�-y���A���m�����#����H˟�U�*ܚ#�4�H�)�f��5!ܪ�d�sco���Euo�o����)�0j�/��
�sD�JV�br���F��𡳤͎b��UQ|d(	���X8�T�ycHn�jۓ�,�p(�+:�[\��4��i�mU4��9R�1o�6Q��*M�D� ���hޥ�P9D�����)r�iBl�Dl�&l�����3��둫?l{J	��mU
�Ȧ�:�;2����Z�?7�is/�߀L�oU�Rh��J�U*�����j���M�ZM��7Cn����٪p���� r�+c�ƴ?�F�vF���f��)\Q��z'-l�6��õ�9$��W���_���2��#�3��m�'Z�h��u�T��T�Q&B��^L�X牖��A<�Pd�,ѝ E��;x�=�����	�G^����zZ@�f�N�;�~�[�X�ky�R�����o�Y/���f�8y(�g��nȭ_�ܥХU�����Ob� �x-ZW����d�]�3�	q7��QS,p�4{��,���wA�����Ytu�5"rW]���[�_?:�ĺ�*�cՉ�Y�F�2�(v<,x��wx��db('��o���s��Z���{bl�i���YK�0Be�ݎ�+�K��:�x�95���
��Ձ��0eb	=2��F$��rŒ��&N)�\��������*��د�4���(�4m��z���ef����m�e�R��.���W�j��.���c���$^�ڜ�{��򉠬N����1Q5e؋]/�>���U�C�k�4��4���i�*��n�H�>g�3��P=.~���r��5�����r&��*��Q��E���f]]z���P�zv:S����p�u�}���i��/�S�]*�*V���~���u�M��c���=��e9Bcdy,.P�bJ�T��#%�������Ͽ���`�i@��.�H����}�Ք56T���ɷ��o�9�u�&6��"�)��oc4dv��Q\U��D_46�V8&8�r�cs��>׻���|e�Y�\�.�?"���/^��%�KTS�}�}n�l,â��������Z�����Ot.�ǻ*�x�̔AfOͱ�Ը�_l��ŧ�����c�����aյ�ۇ؟⡐�#�C%��g]��~S	y�}�� {|Vło��"��t�z��F�u5�|���w#���'�����A{���^s;{�������̑���Ԝ������ Q�'y�Y���eV�R �0(m�}`�����d�HF���(bE�d����wڇ�u,���u�����#��̢\���ߓ�4�M	�c��I��������:��SE;��uJG�tb�d�t�eqi���~y97U:��sW4�F�0��"��='|��0X���%S�2�ijr��6��K�3M%�g�[|�����mA1�����X����1�mq1����Pim�vq�eU�����l[���l�9��kO�Oi��Ϸs����Xo��t��dnD�+��یb�l��佝�k�����/�t0N/
I��$���k���(PI<hvA�"�r�ͧ,X�H��E<[M�غ8�w���^T��-��J��cӆ8�� ��T�#j]�ݕ��øOw���aMc�uD(mdȋ��&+ܥ�R%D^��'F'�2�5V;��~�Z@`c�5M;z��c�1�x�v��QF% �F������+r46W�K].\�� ���n~N����*�x�N�1�����v��O��������v͒���\�oiSF�47]��Ӄ8_���`,\6er��"�.xTӄ����Wv:+Cn�&R��eަZ�x,Y{9�u��,��I�I5�{ի	�+͂fT�_�el�K�Y}�V47HT{�����O�)9r�no`�O{����_�8�\膥G���x� �B=�t7����M�6ƐH"d�f{�"�]1e�"M�6�ov�*�"C��oW�%h���>���O2�^yj\GB�'�<Q�����Y�I�0ם�Ѽ��#��CՕZ+	h���[b��1&͑�y�9	F�9?����<;̎o� �������
qK!�5����i_ʟ]v�ٟG���iXv�ru֥��UIs��d0�;^�4��rj$zP��L&+��+f>��ֺ����̏%I>7jJ��si����s�8�������Y�W���F�'0��~�V����r�gRLO�Q��/��gA��wK	J�L_/3\����L�D��v�GvKĵċ�T��Αg#�k߽{��>����#f�����a!�F�~�i':9�N^��9�(�Đx:�A�^ۆ#>�-�d��g_dR|�n˪�Z��b�l�"�l�Ș0gY��b����lK�YT��@(q
28�&��:�Gw5������@���4��۠��eܫ'|�u��2����\����'�����|�����g~d��y�U)�RC}���uO`I%����FO�t�����LC�׀ ��s]�ZZ�_ψ��^�r�ޏ.�5fJRLU�~z����7�֟޿�F&�sL�
�T�V�Z�&���<�")J�o���}�x�g��}�!YKɘ��|g㨰�<��ܯ!:�5�,;S��wU�g����� BI�n����\�0�
/H��5ǒl����L�9E;պ����K�T�s�Z_=�䨭�$��
�3��`<W�I���_X�Nk=<V��?�Ꭼ����3uMZ�z?�&:�	�߽�5�D��'�&)
�,�_z�C���̇3 a����/���U�T�\�����\�,2[~s�Ǜ�헉��֭������=�8U/���W�ؽ�S��Nu�����t��F�x}�}�(ք�1����
�`��������iw����T�9��j�a6�	"Q������~�v��pK��b§�c��|o�ԽQQN�-�����?ﾔ+$|��E(d-���b���w_�.���c}��]�I�EP���n�/� �e}��	r��%�������=\C5���|e՜?0��3"�����\~��iv��;K]}��2�ϐ�	��?"���-�C�6i�9����h���J��=��,�j��@���Z����m�2ɷ��:�#2�(� �J�պ������u��`9��J�!�N����'�h��}�sO~�8�`�Oit�D�9J�l����ǈ/s^�T����V����V�8,u�4��~p��'�Ξ�[:{OL��'�����1���6��g��~�8l^��K��r�@k�eSүI��+_|u�2��Yʒ�r�qש7	����h����%�.oY��	��?�e1N��-& `��5f�y�t�o��P�7~k� �fv:���ÄO��	���2�z���d��`^�t֏Q6�!���OW��<W�_�A��|���4_>���H�c�cs߁*�����
o�ȥ�z�z?,n~�r@G�����ăW<\�+��d��ُGݝt��"����D��9q��s�>��w͗E�L��/�MQX���H���&Qٕ��n�Jfø���|��ޭ���h��[-�A�����bmk9<K"�~������̕��>zZZ�?���ulnn>6�f�:8{��'��I���mޮf|6�h�lX��f
�tW�o�:
�"Ñn;Ɏ�6΋
?Wx��b=n+�X�ekv?U�_���Nꚤ�}Y}=��ms?^ʘ4��"U~3r��j�&�yv�x�T��c�O,,>|�ƟT�Ԥ�y�^S6�����k{ek�6
vn[󾂪%???�Ivgb��}�4h��I����i>�O����ߋ[(�S��V���亟X�?��v��;[��N�XIS�UV^%������l��6\wװ�--���^�:��o��U.��r�+%,ͤz�bO�-[x,(�]���0��@d��m-b):�� ��̺$��n��c'��ޔ
L�}��S@���(aL�;봡5�]��%��{k�VZ��=R$K���S�VQ�Qv�y�-����'����� "�b���z*���jRI""y>�L�@Ĥ�w��0�#�����˙X��N \�#��vKa�^��6�2�������iwE?�I�s�_7kviU�;�5��6�i�;�a6�ݶ1|0�#�ݽ�'�<|9�J��#){t��uъk���z�H�����G��ms.�Y]�P���X�]E{�'�����&!!�뮍��o�Z�
���j(�{�ۓ[4py�tkk!���SR���}}粳�.�R��ğ��pBh�~��g���%l�������p���v`����Y vtMV�D��v��,¹2o������cB��/�|s�8"�>���hC1a���qPC�Q�ґTv�s1�?>[j�`Y _X��Baĥ���3��W:�����1999]w����ץ��}�.;�K�� ��_��]�뷠8}z��%%��ь����|s}n>�����h���vfɦkZ��}�J`�o���em1b�@X����]�0|��c����٩��[����<����Ȉ/������dz�k�%\br�^�&E�#5��l@�pH��A��5�>���혋��?�4n,������'��>�� '=�<t�����$��C��.�3���՜�A�Њ�G@���/{���&�"$پ��i�o9�UB+'rw�J�5ց�Vsc�?۴�;ءӃ��������8�0T�y1�s�u�tq�o:!����H�#H�)�ĢUJ9@��qV��~���Ç'�,#�ҳ�ez"�y��#����Yzbr��=�y�\����9���c��\��N�A�Bo=x\�b��K}Ü��qb�5��jS�o\���������d��..P���y�� i_io���r����g�����������c�����9���&#.�챜�U4���i�x֜I ��kz�=��;��M��P ��ڳ �-���<��h�������OF�����GTx�B����x�j�f��{��t�+�?�#YE�K>�e����H��Պ:=���=�q�-x��ιa�aP=3�˅W��p�5f��Z���[�FgW�R7x��ۅu����G,n�f�E�����+�	 ��sڗcKO�������u7�:��.�:<C[O�Y&�Kha��T�M&إA�˸�7�����UR6������JB�H�6�(<Xf`�P�$ӺWY���wQ.4����K�;4�/ӿpR~ۏy��#�9��}"f:�oE`<��A�]Ng��Ӌ�h|NL~�ۤk�2񜵅xӥT��xa�B�A�6����S��_�`�'��7̽c�����
�ϷՀ�!�{aj�d��tS���WxS��>@L�캍ݺ�f6�lE 0���V�+m�
���%ҥ�Ů�7Z�T��Ɣ'� 3�X�����u�\ō
-5����:�~ ��~�>Qt\Լ2����������n���$ޝ�g�sbs�>m�
�|��&1w
|Rْd�}� �@G��.�����{`�� R�p�Q��xTB$��dރ�t�(�j	�����QA~~��<��T���ԭ�D�ݽ_d����}_t��d�C�����%�ΕP��䖕'�S�CS���N&S���LjP���&]�nzq�jΐ���X���ޔ1�}���Nd���)u=ԡ�ncS
1��}-��p��;�S'5X�����om�=�޹c��-V�fw�7�,h�}��4d�)���iZ~�e�7�!`rɬ,aׂ�H�&S?֞IpM���l�c-��ÆO$�u�>����I���( �*�{���x���۴VTe��t��M���%k媯�cP(-���J������h�v��\i
�:��;������Ԉ����]0��
%�������_|Y[�T��r!��ҟx�\�І��gZhmܙ;�97�b�;����@2��'�D���+�:�c]o(T�����4���Y��Ϫ�N/rX큄��܌�uTC�c��$R=���YƩ/~�g�}����T�x�\�,��ґ�6y
�&�GO�6��l�*��d�?y�1�忭�<�3\��.�7�A܋֗ڵZ�5�،<[S����1J�Zul1%�rچ:����˯��E�4L}�Zn���8#�z�����~����?l���?������^�}���ND%%���[���s�h}%��1�J'ʉ*��.�F1����d�(E)�ȽjzU��ﵛmdq39`�@�d����x�!ߜ팚��ˤ�@�p�)�l|�rn�w�4�&)H�B�|�7<�̺s�_�Q�r�,�x�D����Ğށ�q�ݲ����K���M~�h��M���3[=��U��Pں�??	=|��B��*��o�3���o�%��SBn\ўLZ��3��D1���Dx�<�p��ԺW v}�ͻ�O6�v.��~~�=�p�ӄ~���iRļk8;;�����'�P�6@k�G�r�i
�HS�yj�(�.��>���m���G��R��F�m!�/��K9-�C�r'����_JP���%)��SO�ҏ�QN���E�Z�
������;�|����,�aʂz�gĥ�W��J�5y@���m����Re
�w���8^M5�p
�,���E��A����ά�{�M"Z�!�+ı7��{�ۋw��O�����n�<m�E���+k���];���lNZHqƋ�;o� [����j@�iց�:�ʠYR�l�4��ZC��9��1�&��2��+v��W��?��:T� ����C�. ���p)��>�>b�����I��ʽ�3�o�|8*��|.81s�^���5{R��5u�/#X�?��ަ���%�Ss���w�z��Thy�����8Fiݔt��3�I��x =���a�ax̒�,1�ݻ��w¹NV��*on\�cb/�i'e�<d��pxG��_����;�{T�;����V��}s�@�2�_,��tvv�-3�F��q<�d�A�m�}5��\�ߣ-�%,)3��W�Ȟ+�U�I��߀V�@PW�*��x���X^�$���;�����/ZR��pCA�BGh�-y>�<��c�*��(*Y�3���}j��#`�2y$&��`�;�>Օ%��#�";�xј�-�%���oMeq��7�"|��	`�c�� ��&�ڶ����:x���}��%ĭx7Wp>[CAם5/�<ڮ�C�U�CC��*tttrQ.���>~����+�J��@�@��f�A��#������\�:��ٙ��]7û*�T��W�>����ggd�!ξc�zc�#�YNV�}�γ"�����	�Ļ�V6q�'��z�`9���l�Y��Sd�L���q����z|�c������0*���纥 �K0�����o��IlY�'W�/��@Z��ȰW�$�V�Z��-6ڔՄ�ݭ�Ȉ"�.��'Fq��1z�u�����ND��`�i�L+�誐�}� ���QΪ�{793\))|���S��ܘ4�n�5�S^
��Q	fۚU�+b4M_;t��߹}q�.���HN���Wy����[9�8��{X�TIF�׾j2Ѫ�ʑ{:�,((�=&���Dgo+�%53�Rs91!�껏�/���j�3w��T�UͶ�%J�9�
G���=[��5rB+r��p�U�>{{��W����R�j3��ۻ��v9��֎/�7�غp�ɫ�?-��b�s����Wm��k	��Y�k��� :�2|9XtB���'��}�������\��)��/�|��Z����}�3i�U�h��2W8��_PT?�'�������6G�a�_yeE�gq/M�N��Yt����w5����])���zW��V�����?gH/�'Q�?e�yr�����?��Әʒ�{%�%��Gh=�W��e���PK   Z�S�Ƽ&�  �     jsons/user_defined.json���o�0�����	��m o��CUm���x�����Y�6��]�߹Y�j�չ���;8�ۣq7H�D���['�J��у�N8��;n��P�����Ň����m7c?)�1���坱;F��<���s�:H�^4%Zu��1,Vʅl0�%�`V�WuJ]�v�ꨥk��c���}T��A�A|��-�HO��rC��ޙ�2�� Ϯͣ?#EV`Q�#��Z&�~LP���nF�����|��U��J�1������ ��u��XH?=k�l����:���'?/��mӻ����
h `B$L��|.h*��&�g_�2��5*����w�/�E/|ɓ\�pTP���$*(�,����FUh yr��U�p�	͓�\�X\�2�)��%IQ�"f���-�p��o�vW�GIn�y\�P��}�����c���?�kiG��M�Jl�N\\���PK
   Z�S$��`�=  �u                  cirkitFile.jsonPK
   L��S1t&�  ב  /             �=  images/3a57aa21-29d3-4406-b48e-ea0158aa2049.pngPK
   Z�S�Ƽ&�  �               �  jsons/user_defined.jsonPK      �   *�    